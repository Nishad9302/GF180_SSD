VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SEVEN_SEG_DECODER
  CLASS BLOCK ;
  FOREIGN SEVEN_SEG_DECODER ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN a
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.840 296.000 22.400 300.000 ;
    END
  END a
  PIN b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 64.400 296.000 64.960 300.000 ;
    END
  END b
  PIN c
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.960 296.000 107.520 300.000 ;
    END
  END c
  PIN d
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 149.520 296.000 150.080 300.000 ;
    END
  END d
  PIN e
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.080 296.000 192.640 300.000 ;
    END
  END e
  PIN f
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.640 296.000 235.200 300.000 ;
    END
  END f
  PIN g
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 277.200 296.000 277.760 300.000 ;
    END
  END g
  PIN i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.520 0.000 38.080 4.000 ;
    END
  END i[0]
  PIN i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 0.000 112.560 4.000 ;
    END
  END i[1]
  PIN i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 186.480 0.000 187.040 4.000 ;
    END
  END i[2]
  PIN i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 0.000 261.520 4.000 ;
    END
  END i[3]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 282.540 ;
      LAYER Metal2 ;
        RECT 21.420 295.700 21.540 296.000 ;
        RECT 22.700 295.700 64.100 296.000 ;
        RECT 65.260 295.700 106.660 296.000 ;
        RECT 107.820 295.700 149.220 296.000 ;
        RECT 150.380 295.700 191.780 296.000 ;
        RECT 192.940 295.700 234.340 296.000 ;
        RECT 235.500 295.700 276.900 296.000 ;
        RECT 21.420 4.300 277.620 295.700 ;
        RECT 21.420 4.000 37.220 4.300 ;
        RECT 38.380 4.000 111.700 4.300 ;
        RECT 112.860 4.000 186.180 4.300 ;
        RECT 187.340 4.000 260.660 4.300 ;
        RECT 261.820 4.000 277.620 4.300 ;
      LAYER Metal3 ;
        RECT 22.330 15.540 274.310 282.380 ;
  END
END SEVEN_SEG_DECODER
END LIBRARY

